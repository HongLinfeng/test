module parity(
    clk,
    rst_n,
    data_in
);
    
endmodule